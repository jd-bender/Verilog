// Jacob Bender
//
// mux4x1.v, 4x1 multiplexor, arrays and composite modules

module DecoderMod(s, o); // module definition
   input [0:1] s;
   output [0:3] o;
   
   wire [0:1] s_inv;
   
   and(o[0], s_inv[1], s_inv[0]);
   and(o[1], s_inv[1], s[0]);
   and(o[2], s[1], s_inv[0]);
   and(o[3], s[1], s[0]);
   not(s_inv[0], s[0]);
   not(s_inv[1], s[1]);
   
endmodule

module MuxMod(s, d, o);
   input [0:1] s;
   input [0:3] d;
   output o;

   wire [0:3] and_out;
   wire [0:3] s_decoded;

   DecoderMod my_decoder(s, s_decoded); // create instance

   and(and_out[0], d[0], s_decoded[0]);
   and(and_out[1], d[1], s_decoded[1]);
   and(and_out[2], d[2], s_decoded[2]);
   and(and_out[3], d[3], s_decoded[3]);
   or(o, and_out[0], and_out[1], and_out[2], and_out[3]);
endmodule

module TestMod;
   reg [0:1] s;
   reg [0:3] d;
   wire o;

   MuxMod my_mux(s, d, o);

   initial begin
      $display("Time\ts[1]\ts[0]\td[0]\td[1]\td[2]\td[3]\to");
      $display("---------------------------------------------------------");
      $monitor("%0d\t%b\t%b\t%b\t%b\t%b\t%b\t%b", $time, s[1], s[0], d[0], d[1], d[2], d[3], o);
   end

   initial begin
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 0; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 0; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 0; d[1] = 1; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 0; d[2] = 1; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 0; d[3] = 1;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 0;
      #1;
      s[1] = 1; s[0] = 1; d[0] = 1; d[1] = 1; d[2] = 1; d[3] = 1;      
      #1; 
   end
endmodule